module frequencyClock(CLOCK_50, pulse);
    input CLOCK_50;
    output pulse;

endmodule