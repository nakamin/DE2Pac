module frequencyLUT(
    input [3:0] note
);
endmodule