module synthesizer(
    input key1_on,
    input [7:0] key1_code,
    input key_2,
    input [7:0] key2_code
);

endmodule