/*
 * map from 8-bit -> 8-bit value for exponential falloff of decay and release
 * in the envelope generator.
 */

 module eight_bit_exponential_decay_lookup (
   input wire [7:0] din,
   output wire [7:0] dout
 );

    assign dout = (
        (din == 8'b00000000) ? 8'hFF : (
        (din == 8'b00000001) ? 8'hF9 : (
        (din == 8'b00000010) ? 8'hF4 : (
        (din == 8'b00000011) ? 8'hEE : (
        (din == 8'b00000100) ? 8'hE9 : (
        (din == 8'b00000101) ? 8'hE4 : (
        (din == 8'b00000110) ? 8'hDF : (
        (din == 8'b00000111) ? 8'hDA : (
        (din == 8'b00001000) ? 8'hD6 : (
        (din == 8'b00001001) ? 8'hD1 : (
        (din == 8'b00001010) ? 8'hCD : (
        (din == 8'b00001011) ? 8'hC8 : (
        (din == 8'b00001100) ? 8'hC4 : (
        (din == 8'b00001101) ? 8'hC0 : (
        (din == 8'b00001110) ? 8'hBB : (
        (din == 8'b00001111) ? 8'hB7 : (
        (din == 8'b00010000) ? 8'hB3 : (
        (din == 8'b00010001) ? 8'hB0 : (
        (din == 8'b00010010) ? 8'hAC : (
        (din == 8'b00010011) ? 8'hA8 : (
        (din == 8'b00010100) ? 8'hA4 : (
        (din == 8'b00010101) ? 8'hA1 : (
        (din == 8'b00010110) ? 8'h9D : (
        (din == 8'b00010111) ? 8'h9A : (
        (din == 8'b00011000) ? 8'h97 : (
        (din == 8'b00011001) ? 8'h93 : (
        (din == 8'b00011010) ? 8'h90 : (
        (din == 8'b00011011) ? 8'h8D : (
        (din == 8'b00011100) ? 8'h8A : (
        (din == 8'b00011101) ? 8'h87 : (
        (din == 8'b00011110) ? 8'h84 : (
        (din == 8'b00011111) ? 8'h81 : (
        (din == 8'b00100000) ? 8'h7E : (
        (din == 8'b00100001) ? 8'h7C : (
        (din == 8'b00100010) ? 8'h79 : (
        (din == 8'b00100011) ? 8'h76 : (
        (din == 8'b00100100) ? 8'h74 : (
        (din == 8'b00100101) ? 8'h71 : (
        (din == 8'b00100110) ? 8'h6F : (
        (din == 8'b00100111) ? 8'h6D : (
        (din == 8'b00101000) ? 8'h6A : (
        (din == 8'b00101001) ? 8'h68 : (
        (din == 8'b00101010) ? 8'h66 : (
        (din == 8'b00101011) ? 8'h63 : (
        (din == 8'b00101100) ? 8'h61 : (
        (din == 8'b00101101) ? 8'h5F : (
        (din == 8'b00101110) ? 8'h5D : (
        (din == 8'b00101111) ? 8'h5B : (
        (din == 8'b00110000) ? 8'h59 : (
        (din == 8'b00110001) ? 8'h57 : (
        (din == 8'b00110010) ? 8'h55 : (
        (din == 8'b00110011) ? 8'h53 : (
        (din == 8'b00110100) ? 8'h52 : (
        (din == 8'b00110101) ? 8'h50 : (
        (din == 8'b00110110) ? 8'h4E : (
        (din == 8'b00110111) ? 8'h4C : (
        (din == 8'b00111000) ? 8'h4B : (
        (din == 8'b00111001) ? 8'h49 : (
        (din == 8'b00111010) ? 8'h48 : (
        (din == 8'b00111011) ? 8'h46 : (
        (din == 8'b00111100) ? 8'h44 : (
        (din == 8'b00111101) ? 8'h43 : (
        (din == 8'b00111110) ? 8'h42 : (
        (din == 8'b00111111) ? 8'h40 : (
        (din == 8'b01000000) ? 8'h3F : (
        (din == 8'b01000001) ? 8'h3D : (
        (din == 8'b01000010) ? 8'h3C : (
        (din == 8'b01000011) ? 8'h3B : (
        (din == 8'b01000100) ? 8'h39 : (
        (din == 8'b01000101) ? 8'h38 : (
        (din == 8'b01000110) ? 8'h37 : (
        (din == 8'b01000111) ? 8'h36 : (
        (din == 8'b01001000) ? 8'h35 : (
        (din == 8'b01001001) ? 8'h33 : (
        (din == 8'b01001010) ? 8'h32 : (
        (din == 8'b01001011) ? 8'h31 : (
        (din == 8'b01001100) ? 8'h30 : (
        (din == 8'b01001101) ? 8'h2F : (
        (din == 8'b01001110) ? 8'h2E : (
        (din == 8'b01001111) ? 8'h2D : (
        (din == 8'b01010000) ? 8'h2C : (
        (din == 8'b01010001) ? 8'h2B : (
        (din == 8'b01010010) ? 8'h2A : (
        (din == 8'b01010011) ? 8'h29 : (
        (din == 8'b01010100) ? 8'h28 : (
        (din == 8'b01010101) ? 8'h28 : (
        (din == 8'b01010110) ? 8'h27 : (
        (din == 8'b01010111) ? 8'h26 : (
        (din == 8'b01011000) ? 8'h25 : (
        (din == 8'b01011001) ? 8'h24 : (
        (din == 8'b01011010) ? 8'h23 : (
        (din == 8'b01011011) ? 8'h23 : (
        (din == 8'b01011100) ? 8'h22 : (
        (din == 8'b01011101) ? 8'h21 : (
        (din == 8'b01011110) ? 8'h20 : (
        (din == 8'b01011111) ? 8'h20 : (
        (din == 8'b01100000) ? 8'h1F : (
        (din == 8'b01100001) ? 8'h1E : (
        (din == 8'b01100010) ? 8'h1E : (
        (din == 8'b01100011) ? 8'h1D : (
        (din == 8'b01100100) ? 8'h1C : (
        (din == 8'b01100101) ? 8'h1C : (
        (din == 8'b01100110) ? 8'h1B : (
        (din == 8'b01100111) ? 8'h1B : (
        (din == 8'b01101000) ? 8'h1A : (
        (din == 8'b01101001) ? 8'h19 : (
        (din == 8'b01101010) ? 8'h19 : (
        (din == 8'b01101011) ? 8'h18 : (
        (din == 8'b01101100) ? 8'h18 : (
        (din == 8'b01101101) ? 8'h17 : (
        (din == 8'b01101110) ? 8'h17 : (
        (din == 8'b01101111) ? 8'h16 : (
        (din == 8'b01110000) ? 8'h16 : (
        (din == 8'b01110001) ? 8'h15 : (
        (din == 8'b01110010) ? 8'h15 : (
        (din == 8'b01110011) ? 8'h14 : (
        (din == 8'b01110100) ? 8'h14 : (
        (din == 8'b01110101) ? 8'h13 : (
        (din == 8'b01110110) ? 8'h13 : (
        (din == 8'b01110111) ? 8'h13 : (
        (din == 8'b01111000) ? 8'h12 : (
        (din == 8'b01111001) ? 8'h12 : (
        (din == 8'b01111010) ? 8'h11 : (
        (din == 8'b01111011) ? 8'h11 : (
        (din == 8'b01111100) ? 8'h11 : (
        (din == 8'b01111101) ? 8'h10 : (
        (din == 8'b01111110) ? 8'h10 : (
        (din == 8'b01111111) ? 8'h10 : (
        (din == 8'b10000000) ? 8'h0F : (
        (din == 8'b10000001) ? 8'h0F : (
        (din == 8'b10000010) ? 8'h0F : (
        (din == 8'b10000011) ? 8'h0E : (
        (din == 8'b10000100) ? 8'h0E : (
        (din == 8'b10000101) ? 8'h0E : (
        (din == 8'b10000110) ? 8'h0D : (
        (din == 8'b10000111) ? 8'h0D : (
        (din == 8'b10001000) ? 8'h0D : (
        (din == 8'b10001001) ? 8'h0C : (
        (din == 8'b10001010) ? 8'h0C : (
        (din == 8'b10001011) ? 8'h0C : (
        (din == 8'b10001100) ? 8'h0C : (
        (din == 8'b10001101) ? 8'h0B : (
        (din == 8'b10001110) ? 8'h0B : (
        (din == 8'b10001111) ? 8'h0B : (
        (din == 8'b10010000) ? 8'h0B : (
        (din == 8'b10010001) ? 8'h0A : (
        (din == 8'b10010010) ? 8'h0A : (
        (din == 8'b10010011) ? 8'h0A : (
        (din == 8'b10010100) ? 8'h0A : (
        (din == 8'b10010101) ? 8'h09 : (
        (din == 8'b10010110) ? 8'h09 : (
        (din == 8'b10010111) ? 8'h09 : (
        (din == 8'b10011000) ? 8'h09 : (
        (din == 8'b10011001) ? 8'h09 : (
        (din == 8'b10011010) ? 8'h08 : (
        (din == 8'b10011011) ? 8'h08 : (
        (din == 8'b10011100) ? 8'h08 : (
        (din == 8'b10011101) ? 8'h08 : (
        (din == 8'b10011110) ? 8'h08 : (
        (din == 8'b10011111) ? 8'h07 : (
        (din == 8'b10100000) ? 8'h07 : (
        (din == 8'b10100001) ? 8'h07 : (
        (din == 8'b10100010) ? 8'h07 : (
        (din == 8'b10100011) ? 8'h07 : (
        (din == 8'b10100100) ? 8'h07 : (
        (din == 8'b10100101) ? 8'h07 : (
        (din == 8'b10100110) ? 8'h06 : (
        (din == 8'b10100111) ? 8'h06 : (
        (din == 8'b10101000) ? 8'h06 : (
        (din == 8'b10101001) ? 8'h06 : (
        (din == 8'b10101010) ? 8'h06 : (
        (din == 8'b10101011) ? 8'h06 : (
        (din == 8'b10101100) ? 8'h06 : (
        (din == 8'b10101101) ? 8'h05 : (
        (din == 8'b10101110) ? 8'h05 : (
        (din == 8'b10101111) ? 8'h05 : (
        (din == 8'b10110000) ? 8'h05 : (
        (din == 8'b10110001) ? 8'h05 : (
        (din == 8'b10110010) ? 8'h05 : (
        (din == 8'b10110011) ? 8'h05 : (
        (din == 8'b10110100) ? 8'h05 : (
        (din == 8'b10110101) ? 8'h04 : (
        (din == 8'b10110110) ? 8'h04 : (
        (din == 8'b10110111) ? 8'h04 : (
        (din == 8'b10111000) ? 8'h04 : (
        (din == 8'b10111001) ? 8'h04 : (
        (din == 8'b10111010) ? 8'h04 : (
        (din == 8'b10111011) ? 8'h04 : (
        (din == 8'b10111100) ? 8'h04 : (
        (din == 8'b10111101) ? 8'h04 : (
        (din == 8'b10111110) ? 8'h04 : (
        (din == 8'b10111111) ? 8'h03 : (
        (din == 8'b11000000) ? 8'h03 : (
        (din == 8'b11000001) ? 8'h03 : (
        (din == 8'b11000010) ? 8'h03 : (
        (din == 8'b11000011) ? 8'h03 : (
        (din == 8'b11000100) ? 8'h03 : (
        (din == 8'b11000101) ? 8'h03 : (
        (din == 8'b11000110) ? 8'h03 : (
        (din == 8'b11000111) ? 8'h03 : (
        (din == 8'b11001000) ? 8'h03 : (
        (din == 8'b11001001) ? 8'h03 : (
        (din == 8'b11001010) ? 8'h03 : (
        (din == 8'b11001011) ? 8'h03 : (
        (din == 8'b11001100) ? 8'h02 : (
        (din == 8'b11001101) ? 8'h02 : (
        (din == 8'b11001110) ? 8'h02 : (
        (din == 8'b11001111) ? 8'h02 : (
        (din == 8'b11010000) ? 8'h02 : (
        (din == 8'b11010001) ? 8'h02 : (
        (din == 8'b11010010) ? 8'h02 : (
        (din == 8'b11010011) ? 8'h02 : (
        (din == 8'b11010100) ? 8'h02 : (
        (din == 8'b11010101) ? 8'h02 : (
        (din == 8'b11010110) ? 8'h02 : (
        (din == 8'b11010111) ? 8'h02 : (
        (din == 8'b11011000) ? 8'h02 : (
        (din == 8'b11011001) ? 8'h02 : (
        (din == 8'b11011010) ? 8'h02 : (
        (din == 8'b11011011) ? 8'h02 : (
        (din == 8'b11011100) ? 8'h02 : (
        (din == 8'b11011101) ? 8'h02 : (
        (din == 8'b11011110) ? 8'h02 : (
        (din == 8'b11011111) ? 8'h01 : (
        (din == 8'b11100000) ? 8'h01 : (
        (din == 8'b11100001) ? 8'h01 : (
        (din == 8'b11100010) ? 8'h01 : (
        (din == 8'b11100011) ? 8'h01 : (
        (din == 8'b11100100) ? 8'h01 : (
        (din == 8'b11100101) ? 8'h01 : (
        (din == 8'b11100110) ? 8'h01 : (
        (din == 8'b11100111) ? 8'h01 : (
        (din == 8'b11101000) ? 8'h01 : (
        (din == 8'b11101001) ? 8'h01 : (
        (din == 8'b11101010) ? 8'h01 : (
        (din == 8'b11101011) ? 8'h01 : (
        (din == 8'b11101100) ? 8'h01 : (
        (din == 8'b11101101) ? 8'h01 : (
        (din == 8'b11101110) ? 8'h01 : (
        (din == 8'b11101111) ? 8'h01 : (
        (din == 8'b11110000) ? 8'h01 : (
        (din == 8'b11110001) ? 8'h01 : (
        (din == 8'b11110010) ? 8'h01 : (
        (din == 8'b11110011) ? 8'h01 : (
        (din == 8'b11110100) ? 8'h01 : (
        (din == 8'b11110101) ? 8'h01 : (
        (din == 8'b11110110) ? 8'h01 : (
        (din == 8'b11110111) ? 8'h01 : (
        (din == 8'b11111000) ? 8'h01 : (
        (din == 8'b11111001) ? 8'h01 : (
        (din == 8'b11111010) ? 8'h01 : (
        (din == 8'b11111011) ? 8'h01 : (
        (din == 8'b11111100) ? 8'h01 : (
        (din == 8'b11111101) ? 8'h01 : (
        (din == 8'b11111110) ? 8'h01 : (
        (din == 8'b11111111) ? 8'h00 : 0
        ))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));

endmodule